//Sam Baker
//10/2023
//Load Store Test

//This is not yet implemented... if that wasnt clear

class load_store_test extends basic_test;








endclass