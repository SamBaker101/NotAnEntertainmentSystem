//Sam Baker
//10/2023
//Basic test to be used with tb_6502_top

//This is not yet implemented... if that wasnt clear

class basic_test;
    


endclass