//Sam Baker
//10/2023
//Basic test to be used with tb_6502_top



class basic_test;
    


endclass