//Sam Baker
//10/2023
//Load Store Test

class load_store_test extends basic_test;








endclass